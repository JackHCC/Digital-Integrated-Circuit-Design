`timescale 1ns  / 10 ps

module carry_out_4 (input  Cin,   input  [3:0] g, p, output Cout);
assign Cout =(( Cin & p[0]&p[1]&p[2]&p[3])     | (g[0]&p[1]&p[2]&p[3])     | (g[1]&p[2]&p[3])      | (g[2]&p[3])       |  g[3] );
endmodule

`timescale 1ns  / 10 ps

module carry_out_16 ( input  Cin,   input  [15:0] g, p, output Cout);
assign Cout = (( Cin &  p[0] &p[1]  &p[2]  &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[0] &p[1]  &p[2]  &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[1] &p[2]  &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[2] &p[3]  &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[3] &p[4]  &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[4] &p[5]  &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[5] &p[6]  &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[6] &p[7]  &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[7] &p[8]  &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[8] &p[9]  &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                       (g[9] &p[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                      (g[10] &p[11] &p[12] &p[13] &p[14] &p[15])  | 
                      (g[11] &p[12] &p[13] &p[14] &p[15])  | 
                      (g[12] &p[13] &p[14] &p[15])  | 
                      (g[13] &p[14] &p[15])  | 
                      (g[14] &p[15])  | 
                      (g[15])
					   );
endmodule
